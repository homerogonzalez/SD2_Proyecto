library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity OR_4 is
    port(OR4_IN: in std_logic_vector(3 downto 0);
            OR4_OUT: out std_logic);
end OR_4;

architecture dataflow of OR_4 is
begin  
    OR4_OUT <= OR4_IN(3) OR OR4_IN(2) OR OR4_IN(1) OR OR4_IN(0);
end dataflow;
            
