module sismin ( 
	a9,
	a8,
	a7,
	a6,
	a5,
	a4,
	a3,
	a2,
	a1,
	a0,
	rw,
	rd,
	wt,
	pe,
	psa,
	psb
	) ;

input  a9;
input  a8;
input  a7;
input  a6;
input  a5;
input  a4;
input  a3;
input  a2;
input  a1;
input  a0;
input  rw;
inout  rd;
inout  wt;
inout  pe;
inout  psa;
inout  psb;
