LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SISMIN IS
PORT(A9,A8,A7,A6,A5,A4,A3,A2,A1,A0,RW: IN STD_LOGIC;
	 RD,WT,PE,PSA,PSB: OUT STD_LOGIC);
END SISMIN;

ARCHITECTURE DATAFLOW OF SISMIN IS
BEGIN

	RD<=NOT RW;

	WT<= RW;

	PE <= NOT (A9 AND A8 AND (NOT A7) AND A6 AND (NOT A5) AND (NOT A4) AND (NOT A3) AND (NOT A2) AND (NOT A1) AND (NOT A0) AND RW);
		--1 1  0 1 0 0  0 0 0 0  0x340

	PSA <= (A9 AND A8 AND (NOT A7) AND (NOT A6) AND A5 AND (NOT A4) AND (NOT A3) AND (NOT A2) AND (NOT A1) AND (NOT A0) AND (NOT RW));
		--1 1  0 0 1 0  0 0 0 0  0x320

	PSB <= (A9 AND A8 AND (NOT A7) AND (NOT A6) AND (NOT A5) AND (NOT A4) AND (NOT A3) AND (NOT A2) AND (NOT A1) AND (NOT A0) AND (NOT RW));
		--1 1  0 0 0 0  0 0 0 0  0x300

END DATAFLOW;
