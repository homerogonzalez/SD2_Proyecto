--alu
